module range

pub struct IntRange {
	start int = 0
	stop int
	step int = 1 

}

pub struct FloatRange {
	start f32 = 1.0
	stop f32
	step f32 = 1.0 

}

pub fn range(range IntRange) []int {
	mut arr := []int{}

	if range.step == 0 {
		eprintln('range: step cannot be zero')
		exit(0)
	}
    if range.start > range.stop {
		if range.step <= -1 {
			for i := range.start; i > range.stop; i += range.step {
			    arr << i
		    }
		}
	}
	for i := range.start; i < range.stop; i += range.step {
		    arr << i
	}
	return arr
}

pub fn range_float(float FloatRange) []f32 {
	mut arr := []f32{}

	if float.step == 0 {
		eprintln('range: step cannot be zero')
		exit(0)
	}
    if float.start > float.stop {
			for i := float.start; i > float.stop; i += float.step {
			    arr << i
		    }
	}
	for i := float.start; i < float.stop; i += float.step {
		    arr << i
	}
	return arr
}
